TACS (PSpice format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             ** 
**      (c) DesignSoft, Inc.        **          
**     www.designsoftware.com       **
**************************************
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\EXAMPLES\SPICE\TSPICE.LIB"
.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\Operational Amplifiers.LIB"
.LIB
.TEMP 27
.AC DEC 20 10 1MEG
.TRAN 200U 100M UIC
.DC LIN VG1 0 1 10M

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE I(VAM1) V([VF2])

VG1         3 228 DC 0 AC 1 0
+ SIN( 0 1.5 80 0 0 0 )
VG1_DC      228 4 3.5
VAM1        20 VF2 ; AmperMeter
VS2         0 4 36
VS1         22 0 36
XU1         1 2 LM4040_NA5P0_0
+ PARAMS: TOL=0
XU4         5 6 LM4040_NA10P0_0
+ PARAMS: TOL=0
XU12        5 7 LM4040_NA2P5_0
+ PARAMS: TOL=0
XU9         8 4 LM4040_NA10P0_0
+ PARAMS: TOL=0
XU6         7 9 5 11 10 TLC2252_0
DLED2       12 4  D_CQX35A_1 
XU7         3 13 1 4 14 TLC2252_0
DLED1       15 16  D_CQX35A_1 
XU8         3 17 1 4 18 TLC2252_0
XU2         11 7 5 7 19 TLC2252_0
C2          4 1 1U 
R16         12 22 75K 
R15         23 22 75K 
R14         15 23 75K 
R13         24 14 75K 
R12         4 24 75K 
R11         8 0 36K 
R10         0 6 36K 
R9          11 7 7.15K 
R8          9 5 1K 
C1          4 2 1U 
R7          4 13 7.15K 
R6          13 2 75K 
R5          25 4 86.6 
R4          17 25 1K 
R3          26 27 2.2K 
R2          20 26 2.2K 
R1          0 VF2 4K 
QT6         27 10 9  Q__PNP_P_1 
QT5         27 18 17  Q__NPN_N_1 
QT4         16 24 4  Q__NPN_N_1 
QT3         0 6 11  Q__PNP_P_1 
QT2         5 23 22  Q__PNP_P_1 
QT1         0 8 1  Q__NPN_N_1 

.MODEL D_CQX35A_1 D( IS=5.62P N=2.8 BV=5 IBV=100U RS=420M 
+      CJO=35P VJ=750M M=330M FC=500M TT=100N 
+      EG=1.11 XTI=3 KF=0 AF=1 )
.MODEL Q__PNP_P_1 PNP( IS=9.85F NF=1 NR=1 RE=3.18 RC=1 
+      RB=10 VAF= 1.00000000000000E+0030 VAR= 1.00000000000000E+0030 ISE=0 ISC=0 
+      ISS=0 NE=1.5 NC=1.5 NS=1 BF=567 
+      BR=5 IKF=0 IKR=0 CJC=8.96P CJE=9.35P 
+      CJS=0 VJC=615M VJE=991M VJS=750M MJC=330M 
+      MJE=426M MJS=0 TF=531P TR=69N EG=1.11 
+      KF=0 AF=1 )
.MODEL Q__NPN_N_1 NPN( IS=12.6F NF=991M NR=991M RE=305M RC=1 
+      RB=10 VAF= 1.00000000000000E+0030 VAR= 1.00000000000000E+0030 ISE=0 ISC=0 
+      ISS=0 NE=1.5 NC=1.5 NS=1 BF=100 
+      BR=5 IKF=0 IKR=0 CJC=10.4P CJE=14.8P 
+      CJS=0 VJC=100M VJE=100M VJS=750M MJC=278M 
+      MJE=237M MJS=0 TF=531P TR=69N EG=1.11 
+      KF=0 AF=1 )

* PSPICE MODEL EDITOR - VERSION 16.0.0
*$
*LM4040_N
*****************************************************************************
*  (C) COPYRIGHT 2013 TEXAS INSTRUMENTS INCORPORATED. ALL RIGHTS RESERVED.
*****************************************************************************
** THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.
** TI AND ITS LICENSORS AND SUPPLIERS MAKE NO WARRANTIES, EITHER EXPRESSED
** OR IMPLIED, WITH RESPECT TO THIS MODEL, INCLUDING THE WARRANTIES OF 
** MERCHANTABILITY OR FITNESS FOR A PARTICULAR PURPOSE. THE MODEL IS
** PROVIDED SOLELY ON AN "AS IS" BASIS. THE ENTIRE RISK AS TO ITS QUALITY
** AND PERFORMANCE IS WITH THE CUSTOMER.
*****************************************************************************
*
** RELEASED BY: WEBENCH DESIGN CENTER,TEXAS INSTRUMENTS INC.
* PART: LM4040_N
* DATE: 10APR2013
* MODEL TYPE: TRANSIENT
* SIMULATOR: PSPICE
* SIMULATOR VERSION: 16.0.0
* EVM ORDER NUMBER: N/A
* EVM USERS GUIDE: N/A
* DATASHEET: SNOS633G�MAY 2004�REVISED JULY 2012
*
* MODEL VERSION: FINAL 1.00
*
*****************************************************************************
*
* UPDATES:
*
* FINAL 1.00
* RELEASE TO WEB.
*
******************************************************************************
.SUBCKT LM4040_NA5P0_0  V+ V-  PARAMS: TOL=0
C_CSTART         V- START  400NF  TC=0,0 
Q_Q22         N03098 N01931 V- NPN1X 
Q_Q7         N02184 VC_Q2 N01786 NPN1X 
Q_Q12         N02229 N03098 N04190 NPN1X 
Q_Q13         N04160 N04160 N04190 NPN1X 10
Q_Q3         VC_Q3 VB_Q3 VE NPN1X 10
Q_Q5         VC_Q3 N01129 N01136 PNPL1X 1.8
Q_Q6         N01129 N01129 N01136 PNPL1X 1.8
C_C3         N03098 N01136  3PF  TC=0,0 
Q_Q23         N01136 N01136 N08107 NPN1X 
R_R10         N01129 N01786  60K TC=0,0 
Q_Q15         N04160 N02229 N01136 PNPL1X 10
R_R1TOR5         N07686 N01136  30.5K TC=0,0 
R_R15         N01931 Q20B  66K TC=0,0 
Q_Q14         N02229 N02229 N01136 PNPL1X 1
Q_Q20         N01533 Q20B V- NPN1X 
R_R6         VB_Q2 N07686  20K TC=0,0 
C_CX         V- N01136  1PF  TC=0,0 
C_C2         VC_Q3 N02514  6PF  TC=0,0 
E_ESTART         N30465 V- VALUE { MAX(0.4*(1-V(VB_Q2, VB_Q3)/.05), 0)+V(Q20B)
+  }
Q_Q1         V- FB_TEMP Q1E PNPV1X 5
Q_Q17         N01533 FB_TEMP Q1E PNPL1X 1
R_RX6         V+ N01136  1000 TC=0,0 
Q_Q19         Q20B VE N08426 PNPL1X 1
R_R8         Q1E VB_Q3  45K TC=0,0 
Q_Q16         N01136 N04160 V- NPN1X 10
Q_Q4         VC_Q2 N01129 N01136 PNPL1X 1.8
R_R13         Q20B N01533  40K TC=0,0 
R_RSTART0         START N30465  200 TC=0,0 
R_R11         N02514 N02184  100K TC=0,0 
R_R14         N01755 V-  3.3K TC=0,0 
Q_Q11         N03098 N02514 N01136 PNPL1X 1.8
Q_Q21         N01786 Q20B N01755 NPN1X 6.75
Q_Q24         N01136 N07686 N08116 NPN1X 
Q_Q8         N02514 VC_Q3 N01786 NPN1X 
Q_Q2         VC_Q2 VB_Q2 VE NPN1X 
Q_Q10         N02514 N02184 N01136 PNPL1X 3.1
Q_Q9         N02184 N02184 N01136 PNPL1X 3.1
R_R18         Q1E N08116  69K TC=0,0 
R_R59         N01136 N08426  51K TC=0,0 
R_R12         N01505 V-  6K TC=0,0 
L_LX1         N01136 V+  10UH  
R_R16         N04190 V-  1K TC=0,0 
Q_Q18         VE Q20B N01505 NPN1X 
R_RSTART1         Q20B START  20K TC=0,0 
R_R17         N08116 N08107  130K TC=0,0 
R_R7         VB_Q3 VB_Q2  10K TC=0,0 
C_C1         VC_Q2 N03098  3PF  TC=0,0 
R_R19       V+ FB_TEMP    {IF({TOL}==0,162218.6,IF({TOL}>0,162065.9, 162371.3 ))} 
R_R20       FB_TEMP V-  500K 
.MODEL NPN1X NPN IS=13.84E-18 BF=130 TR=8NS
.MODEL PNPV1X PNP IS=261.8E-18 BF=222
.MODEL PNPL1X PNP  IS=48E-18 BF=63
.MODEL MENABLE NMOS LEVEL 1
+ VTO 0
+ KP 20.000000E-06
+ PHI 0.6
+ IS 10.000000E-15
+ PB     .8          
+ PBSW     .8          
+ UCRIT   10.000000E+03 
+ DIOMOD    1             
*+ VDD    5            
*+ XPART    0            
*
*
.MODEL DIDEAL D IS=0.001P N=0.01 RS=0 IKF=0 XTI=2 EG=1.11 CJO=0
+               M=0.33 VJ=1 FC=0.5 ISR=0.1N NR=2 BV=75 IBV=1E-10 TT=0
*
*
.ENDS LM4040_NA5P0_0 
*$


* PSPICE MODEL EDITOR - VERSION 16.0.0
*$
*LM4040_N
*****************************************************************************
*  (C) COPYRIGHT 2013 TEXAS INSTRUMENTS INCORPORATED. ALL RIGHTS RESERVED.
*****************************************************************************
** THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.
** TI AND ITS LICENSORS AND SUPPLIERS MAKE NO WARRANTIES, EITHER EXPRESSED
** OR IMPLIED, WITH RESPECT TO THIS MODEL, INCLUDING THE WARRANTIES OF 
** MERCHANTABILITY OR FITNESS FOR A PARTICULAR PURPOSE. THE MODEL IS
** PROVIDED SOLELY ON AN "AS IS" BASIS. THE ENTIRE RISK AS TO ITS QUALITY
** AND PERFORMANCE IS WITH THE CUSTOMER.
*****************************************************************************
*
** RELEASED BY: WEBENCH DESIGN CENTER,TEXAS INSTRUMENTS INC.
* PART: LM4040_N
* DATE: 10APR2013
* MODEL TYPE: TRANSIENT
* SIMULATOR: PSPICE
* SIMULATOR VERSION: 16.0.0
* EVM ORDER NUMBER: N/A
* EVM USERS GUIDE: N/A
* DATASHEET: SNOS633G�MAY 2004�REVISED JULY 2012
*
* MODEL VERSION: FINAL 1.00
*
*****************************************************************************
*
* UPDATES:
*
* FINAL 1.00
* RELEASE TO WEB.
*
******************************************************************************
.SUBCKT LM4040_NA10P0_0   V+ V- PARAMS: TOL=0
C_CSTART         V- START  400NF  TC=0,0 
Q_Q22         N03098 N01931 V- NPN1X 
Q_Q7         N02184 VC_Q2 N01786 NPN1X 
Q_Q12         N02229 N03098 N04190 NPN1X 
Q_Q13         N04160 N04160 N04190 NPN1X 10
Q_Q3         VC_Q3 VB_Q3 VE NPN1X 10
Q_Q5         VC_Q3 N01129 N01136 PNPL1X 1.8
Q_Q6         N01129 N01129 N01136 PNPL1X 1.8
C_C3         N03098 N01136  3PF  TC=0,0 
Q_Q23         N01136 N01136 N08107 NPN1X 
R_R10         N01129 N01786  60K TC=0,0 
Q_Q15         N04160 N02229 N01136 PNPL1X 10
R_R1TOR5         N07686 N01136  30.5K TC=0,0 
R_R15         N01931 Q20B  66K TC=0,0 
Q_Q14         N02229 N02229 N01136 PNPL1X 1
Q_Q20         N01533 Q20B V- NPN1X 
R_R6         VB_Q2 N07686  20K TC=0,0 
C_CX         V- N01136  1PF  TC=0,0 
C_C2         VC_Q3 N02514  6PF  TC=0,0 
E_ESTART         N30465 V- VALUE { MAX(0.4*(1-V(VB_Q2, VB_Q3)/.05), 0)+V(Q20B)
+  }
Q_Q1         V- FB_TEMP Q1E PNPV1X 5
Q_Q17         N01533 FB_TEMP Q1E PNPL1X 1
R_RX6         V+ N01136  1000 TC=0,0 
Q_Q19         Q20B VE N08426 PNPL1X 1
R_R8         Q1E VB_Q3  45K TC=0,0 
Q_Q16         N01136 N04160 V- NPN1X 10
Q_Q4         VC_Q2 N01129 N01136 PNPL1X 1.8
R_R13         Q20B N01533  40K TC=0,0 
R_RSTART0         START N30465  225 TC=0,0 
R_R11         N02514 N02184  100K TC=0,0 
R_R14         N01755 V-  3.3K TC=0,0 
Q_Q11         N03098 N02514 N01136 PNPL1X 1.8
Q_Q21         N01786 Q20B N01755 NPN1X 6.75
Q_Q24         N01136 N07686 N08116 NPN1X 
Q_Q8         N02514 VC_Q3 N01786 NPN1X 
Q_Q2         VC_Q2 VB_Q2 VE NPN1X 
Q_Q10         N02514 N02184 N01136 PNPL1X 3.1
Q_Q9         N02184 N02184 N01136 PNPL1X 3.1
R_R18         Q1E N08116  69K TC=0,0 
R_R59         N01136 N08426  51K TC=0,0 
R_R12         N01505 V-  6K TC=0,0 
L_LX1         N01136 V+  10UH  
R_R16         N04190 V-  1K TC=0,0 
Q_Q18         VE Q20B N01505 NPN1X 
R_RSTART1         Q20B START  20K TC=0,0 
R_R17         N08116 N08107  130K TC=0,0 
R_R7         VB_Q3 VB_Q2  10K TC=0,0 
C_C1         VC_Q2 N03098  3PF  TC=0,0 
R_R19       V+ FB_TEMP {IF({TOL}==0,111529.8505,IF({TOL}>0,111504.701,111555))} 
R_R20       FB_TEMP V-  800K
.MODEL NPN1X NPN IS=13.84E-18 BF=130 TR=8NS
.MODEL PNPV1X PNP IS=261.8E-18 BF=222
.MODEL PNPL1X PNP  IS=48E-18 BF=63
.MODEL MENABLE NMOS LEVEL 1
+ VTO 0
+ KP 20.000000E-06
+ PHI 0.6
+ IS 10.000000E-15
+ PB     .8          
+ PBSW     .8          
+ UCRIT   10.000000E+03 
+ DIOMOD    1             
*+ VDD    5            
*+ XPART    0            
*
*
.MODEL DIDEAL D IS=0.001P N=0.01 RS=0 IKF=0 XTI=2 EG=1.11 CJO=0
+               M=0.33 VJ=1 FC=0.5 ISR=0.1N NR=2 BV=75 IBV=1E-10 TT=0
*
*
.ENDS  LM4040_NA10P0_0 
*$


* PSPICE MODEL EDITOR - VERSION 16.0.0
*$
*LM4040_N
*****************************************************************************
*  (C) COPYRIGHT 2013 TEXAS INSTRUMENTS INCORPORATED. ALL RIGHTS RESERVED.
*****************************************************************************
** THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.
** TI AND ITS LICENSORS AND SUPPLIERS MAKE NO WARRANTIES, EITHER EXPRESSED
** OR IMPLIED, WITH RESPECT TO THIS MODEL, INCLUDING THE WARRANTIES OF 
** MERCHANTABILITY OR FITNESS FOR A PARTICULAR PURPOSE.  THE MODEL IS
** PROVIDED SOLELY ON AN "AS IS" BASIS.  THE ENTIRE RISK AS TO ITS QUALITY
** AND PERFORMANCE IS WITH THE CUSTOMER
*****************************************************************************
*
** RELEASED BY: WEBENCH DESIGN CENTER,TEXAS INSTRUMENTS INC.
* PART: LM4040_N
* DATE: 10APR2013
* MODEL TYPE: TRANSIENT
* SIMULATOR: PSPICE
* SIMULATOR VERSION: 16.0.0
* EVM ORDER NUMBER: N/A
* EVM USERS GUIDE: N/A
* DATASHEET: SNOS633G�MAY 2004�REVISED JULY 2012
*
* MODEL VERSION: FINAL 1.00
*
*****************************************************************************
*
* UPDATES:
*
* FINAL 1.00
* RELEASE TO WEB.
*
******************************************************************************
.SUBCKT LM4040_NA2P5_0   V+ V- PARAMS: TOL=0
C_CSTART         V- START   100NF  TC=0,0 
Q_Q22         N03098 N01931 V- NPN1X 
Q_Q7         N02184 VC_Q2 N01786 NPN1X 
Q_Q12         N02229 N03098 N04190 NPN1X 
Q_Q13         N04160 N04160 N04190 NPN1X 10
Q_Q3         VC_Q3 VB_Q3 VE NPN1X 10
Q_Q5         VC_Q3 N01129 N01136 PNPL1X 1.8
Q_Q6         N01129 N01129 N01136 PNPL1X 1.8
C_C3         N03098 N01136  3PF  TC=0,0 
Q_Q23         N01136 N01136 N08107 NPN1X 
R_R10         N01129 N01786  60K TC=0,0 
Q_Q15         N04160 N02229 N01136 PNPL1X 10
R_R1TOR5         N07686 N01136  30.5K TC=0,0 
R_R15         N01931 Q20B  66K TC=0,0 
Q_Q14         N02229 N02229 N01136 PNPL1X 1
Q_Q20         N01533 Q20B V- NPN1X 
R_R6         VB_Q2 N07686  20K TC=0,0 
C_CX         V- N01136  1PF  TC=0,0 
C_C2         VC_Q3 N02514  6PF  TC=0,0 
E_ESTART         N30465 V- VALUE { MAX(0.4*(1-V(VB_Q2, VB_Q3)/.05), 0)+V(Q20B)
+  }
Q_Q1         V- FB_TEMP Q1E PNPV1X 5
Q_Q17         N01533 FB_TEMP Q1E PNPL1X 1
R_RX6         V+ N01136  1000 TC=0,0 
Q_Q19         Q20B VE N08426 PNPL1X 1
R_R8         Q1E VB_Q3  45K TC=0,0 
Q_Q16         N01136 N04160 V- NPN1X 10
Q_Q4         VC_Q2 N01129 N01136 PNPL1X 1.8
R_R13         Q20B N01533  40K TC=0,0 
R_RSTART0         START N30465 180 TC=0,0 
R_R11         N02514 N02184  100K TC=0,0 
R_R14         N01755 V-  3.3K TC=0,0 
Q_Q11         N03098 N02514 N01136 PNPL1X 1.8
Q_Q21         N01786 Q20B N01755 NPN1X 6.75
Q_Q24         N01136 N07686 N08116 NPN1X 
Q_Q8         N02514 VC_Q3 N01786 NPN1X 
Q_Q2         VC_Q2 VB_Q2 VE NPN1X 
Q_Q10         N02514 N02184 N01136 PNPL1X 3.1
Q_Q9         N02184 N02184 N01136 PNPL1X 3.1
R_R18         Q1E N08116  69K TC=0,0 
R_R59         N01136 N08426  51K TC=0,0 
R_R12         N01505 V-  6K TC=0,0 
L_LX1         N01136 V+  10UH  
R_R16         N04190 V-  1K TC=0,0 
Q_Q18         VE Q20B N01505 NPN1X 
R_RSTART1         Q20B START  20K TC=0,0 
R_R17         N08116 N08107  130K TC=0,0 
R_R7         VB_Q3 VB_Q2  10K TC=0,0 
C_C1         VC_Q2 N03098  3PF  TC=0,0 
R_R19       V+ FB_TEMP  {IF({TOL}==0,483.14225K,IF({TOL}>0,4.826578E5,4.836267E5))}
R_R20       FB_TEMP V-  500K
.MODEL NPN1X NPN IS=13.84E-18 BF=130 TR=8NS
.MODEL PNPV1X PNP IS=261.8E-18 BF=222
.MODEL PNPL1X PNP  IS=48E-18 BF=63
.MODEL MENABLE NMOS LEVEL 1
+ VTO 0
+ KP 20.000000E-06
+ PHI 0.6
+ IS 10.000000E-15
+ PB     .8          
+ PBSW     .8          
+ UCRIT   10.000000E+03 
+ DIOMOD    1             
*+ VDD    5            
*+ XPART    0            
*
*
.MODEL DIDEAL D IS=0.001P N=0.01 RS=0 IKF=0 XTI=2 EG=1.11 CJO=0
+               M=0.33 VJ=1 FC=0.5 ISR=0.1N NR=2 BV=75 IBV=1E-10 TT=0
*
*
.ENDS  LM4040_NA2P5_0 
*$


.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\Operational Amplifiers.LIB"
* TLC2252 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 01/12/95 AT 08:26
* REV (N/A) (10V MODEL) (LEVEL II)
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC2252_0   1 2 3 4 5
*
C1   11 12 6.043E-12
C2    6  7 50.00E-12
CPSR 85 86 7.96E-9
DCM+ 81 82 DX
DCM- 83 81 DX
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
ECMR 84 99 (2,99) 1
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
EPSR 85 0 POLY(1) (3,4) -1736E-6  173.6E-6
ENSE 89 2 POLY(1) (88,0) 200E-6  1
FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 200E6 -30E6 30E6 30E6 -30E6 30E6
GA    6  0 11 12 28.27E-6
GCM 0  6 10 99 2.635E-9
GPSR 85 86 (85,86) 100E-6
GRD1 60 11 (60,11) 28.273E-6
GRD2 60 12 (60,12) 28.273E-6
HLIM 90 0 VLIM 1K
HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
IRP 3 4 34E-6
ISS   3 10 DC 6.000E-6
IIO 2 0 .5E-12
I1 88 0 1E-21
J1   11  89 10 JX
J2   12  80 10 JX
R2    6  9 100.0E3
RCM 84 81 1K
RN1 88 0 100
RO1   8  5 70
RO2   7 99 50
RSS  10 99 33.33E6
VAD 60 4 -.5
VCM+ 82 99 3.6
VCM- 83 99 -4.7
VB    9  0 DC 0
VC 3 53 DC .656
VE   54  4 DC .656
VLIM  7  8 DC 0
VLP  91  0 DC -.234
VLN 0 92 DC 7.5
VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=500.0E-15 BETA=360E-6 VTO=-.023 KF=8.6E-18)
.ENDS


.END
